`ifndef ALU4_DEFINES_SVH
`define ALU4_DEFINES_SVH

`define ALU_OP_ADD  3'b000
`define ALU_OP_SUB  3'b001
`define ALU_OP_AND  3'b010
`define ALU_OP_OR   3'b011
`define ALU_OP_XOR  3'b100

`endif
